(* blackbox *)
module bufgctrl(i, s, ce, ignore, o);
input [1:0] i;
input [1:0] s;
input [1:0] ce;
input [1:0] ignore;
output o;
endmodule

