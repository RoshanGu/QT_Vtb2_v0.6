(* blackbox *)
module xadder(a_xor_b, a_and_b, cin, cout, sumout);
input a_xor_b, a_and_b, cin;
output cout, sumout;
endmodule
