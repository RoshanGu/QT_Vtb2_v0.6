module lut8(A6_1, B6_1, C6_1, D6_1, AX, BX, CX, F8);
input [5:0] A6_1;
input [5:0] B6_1;
input [5:0] C6_1;
input [5:0] D6_1;
input AX, BX, CX;
output F8;
endmodule


