module lut7(A6_1, B6_1, AX, F7);
input [5:0] A6_1;
input [5:0] B6_1;
input AX;
output F7;
endmodule
